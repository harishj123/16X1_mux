interface mux_16x1_interface(input logic clk);
  logic rst;
  logic [15:0] [31:0] i;
  logic [3:0] s;
  logic [31:0] y;
endinterface
